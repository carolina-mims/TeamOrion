`timescale 1 ns/100 ps
module testbench_GameController( );

    reg Passed_s, LoadPlayerIn_s, GameStartButton_s, Clk_s, Rst_s, TimerTimeout_s, FinGen_s, TwoSecTimeout_s;
    reg [3:0] PlayerNum_s;
    reg [3:0] RAMOutput_s;
    reg [4:0] PlayerID_s;
    wire TimerReconfig_s, TimerEnable_s, GoGen_s, TwoSecEnable_s;
    wire [3:0] Diff_s;
    wire [4:0] SeqAddr_s;
    wire [3:0] DispDigit_s;
    wire Logout_s;
    wire PersonalWin_s, GlobalWinner_s;

    always
      begin
        Clk_s = 1'b0;
        #10;
        Clk_s = 1'b1;
        #10;
      end

    GameController DUT_GameController(Passed_s, LoadPlayerIn_s, GameStartButton_s, Clk_s, Rst_s, TimerReconfig_s, TimerEnable_s, TimerTimeout_s, GoGen_s, FinGen_s, SeqAddr_s, Diff_s, PlayerNum_s, RAMOutput_s, DispDigit_s, TwoSecEnable_s, TwoSecTimeout_s, PlayerID_s, PersonalWin_s, GlobalWinner_s, Logout_s);

    initial
      begin
        Passed_s = 1'b0;
        LoadPlayerIn_s = 1'b0;
        GameStartButton_s = 1'b0;
        Rst_s = 1'b1;
        TimerTimeout_s = 1'b0;
        FinGen_s = 1'b0;
        TwoSecTimeout_s = 1'b0;
        PlayerNum_s = 4'b0000;
        RAMOutput_s = 4'b1111;
        PlayerID_s = 5'b00000;
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 Rst_s = 1'b0;

        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 Rst_s = 1'b1;
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 Passed_s = 1'b1;
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 PlayerNum_s = 4'b0001;
        GameStartButton_s = 4'b0001;
        @(posedge Clk_s);
        #5 GameStartButton_s = 4'b0000;
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 GameStartButton_s = 4'b0001;
        @(posedge Clk_s);
        #5 GameStartButton_s = 4'b0000;
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 FinGen_s = 1'b1;
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 GameStartButton_s = 4'b0001;
        @(posedge Clk_s);
        #5 GameStartButton_s = 4'b0000;
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 RAMOutput_s = 4'b1001;
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 TwoSecTimeout_s = 1'b1;
        @(posedge Clk_s);
        #5 TwoSecTimeout_s = 1'b0;
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 RAMOutput_s = 4'b1001;
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 TwoSecTimeout_s = 1'b1;
        @(posedge Clk_s);
        #5 TwoSecTimeout_s = 1'b0;
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 RAMOutput_s = 4'b1011;
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 TwoSecTimeout_s = 1'b1;
        @(posedge Clk_s);
        #5 TwoSecTimeout_s = 1'b0;
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 RAMOutput_s = 4'b1101;
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 TwoSecTimeout_s = 1'b1;
        @(posedge Clk_s);
        #5 TwoSecTimeout_s = 1'b0;
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 TwoSecTimeout_s = 1'b1;
        @(posedge Clk_s);
        #5 TwoSecTimeout_s = 1'b0;
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 GameStartButton_s = 4'b0001;
        @(posedge Clk_s);
        #5 GameStartButton_s = 4'b0000;
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 RAMOutput_s = 4'b1001;
        PlayerNum_s = 4'b1001;
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 LoadPlayerIn_s = 4'b0001;
        @(posedge Clk_s);
        #5 LoadPlayerIn_s = 4'b0000;
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 RAMOutput_s = 4'b1011;
        PlayerNum_s = 4'b1001;
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 LoadPlayerIn_s = 4'b0001;
        @(posedge Clk_s);
        #5 LoadPlayerIn_s = 4'b0000;
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        #5 TimerTimeout_s = 4'b0001;
        @(posedge Clk_s);
        #5 TimerTimeout_s = 4'b0000;
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
        @(posedge Clk_s);
  end

endmodule
